`timescale 1ns / 1ps

module ascii_rom2(
input clk,
input wire [5:0] letterNum,
input wire [3:0] row,
output reg [7:0]data
    );
    
    (*rom_style = "block" *)
    
    always @ (*)
        case(letterNum)
        6'b000000: begin //L
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b00000000;	//
                4'h3: data = 8'b00000000;	//
                4'h4: data = 8'b00000000;	//
                4'h5: data = 8'b00000000;	//
                4'h6: data = 8'b00000000;	//
                4'h7: data = 8'b00000000;	//
                4'h8: data = 8'b00000000;	//
                4'h9: data = 8'b00000000;	//
                4'ha: data = 8'b00000000;	//
                4'hb: data = 8'b00000000;	//
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b000001: begin //A
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b00010000;	//   *
                4'h3: data = 8'b00111000;	//  ***
                4'h4: data = 8'b01101100;	// ** **   
                4'h5: data = 8'b11000110;	//**   **   
                4'h6: data = 8'b11000110;	//**   **
                4'h7: data = 8'b11111110;	//*******
                4'h8: data = 8'b11111110;	//*******
                4'h9: data = 8'b11000110;	//**   **
                4'ha: data = 8'b11000110;	//**   **
                4'hb: data = 8'b11000110;	//**   **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
             endcase
        end
        6'b000010: begin //B
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111100;	//******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **   
                4'h6: data = 8'b11111100;	//******
                4'h7: data = 8'b11111100;	//******
                4'h8: data = 8'b11000110;	//**   **
                4'h9: data = 8'b11000110;	//**   **
                4'ha: data = 8'b11111110;	//*******
                4'hb: data = 8'b11111100;	//******
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b000011: begin // C
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b01111100;	// *****
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000000;	//**
                4'h5: data = 8'b11000000;	//**   
                4'h6: data = 8'b11000000;	//**
                4'h7: data = 8'b11000000;	//**
                4'h8: data = 8'b11000000;	//** 
                4'h9: data = 8'b11000000;	//** 
                4'ha: data = 8'b11111110;	//*******
                4'hb: data = 8'b01111100;	// *****
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;    //
                endcase
        end
        6'b000100: begin //D
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111100;	//******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **   
                4'h6: data = 8'b11000110;	//**   **
                4'h7: data = 8'b11000110;	//**   **
                4'h8: data = 8'b11000110;	//**   ** 
                4'h9: data = 8'b11000110;	//**   ** 
                4'ha: data = 8'b11111110;	//*******
                4'hb: data = 8'b11111100;	//******
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b000101: begin //E
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111110;	//*******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000000;	//**
                4'h5: data = 8'b11000000;	//**   
                4'h6: data = 8'b11111100;	//******
                4'h7: data = 8'b11111100;	//******
                4'h8: data = 8'b11000000;	//** 
                4'h9: data = 8'b11000000;	//** 
                4'ha: data = 8'b11111110;	//*******
                4'hb: data = 8'b11111110;	//*******
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b000110: begin //F
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111110;	//*******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000000;	//**
                4'h5: data = 8'b11000000;	//**   
                4'h6: data = 8'b11111100;	//******
                4'h7: data = 8'b11111100;	//******
                4'h8: data = 8'b11000000;	//** 
                4'h9: data = 8'b11000000;	//** 
                4'ha: data = 8'b11000000;	//**
                4'hb: data = 8'b11000000;	//**
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b000111: begin //G
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b01111100;	// *****
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000000;	//**
                4'h5: data = 8'b11000000;	//**   
                4'h6: data = 8'b11111110;	//*******
                4'h7: data = 8'b11111110;	//*******
                4'h8: data = 8'b11000110;	//**   **
                4'h9: data = 8'b11000110;	//**   **
                4'ha: data = 8'b11111110;	//*******
                4'hb: data = 8'b01111110;	// ******
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b001000: begin //H
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000110;	//**   **
                4'h3: data = 8'b11000110;	//**   **
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **
                4'h6: data = 8'b11111110;	//*******
                4'h7: data = 8'b11111110;	//*******
                4'h8: data = 8'b11000110;	//**   **
                4'h9: data = 8'b11000110;	//**   **
                4'ha: data = 8'b11000110;	//**   **
                4'hb: data = 8'b11000110;	//**   **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//  
                endcase
        end
        6'b001001: begin //I
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111110;	//*******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b00110000;	//  **
                4'h5: data = 8'b00110000;	//  **
                4'h6: data = 8'b00110000;	//  **
                4'h7: data = 8'b00110000;	//  **
                4'h8: data = 8'b00110000;	//  **
                4'h9: data = 8'b00110000;	//  **
                4'ha: data = 8'b11111110;	//*******
                4'hb: data = 8'b11111110;	//*******
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b001010: begin //J
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111110;	//*******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b00011000;	//   **
                4'h5: data = 8'b00011000;	//   **
                4'h6: data = 8'b00011000;	//   **
                4'h7: data = 8'b00011000;	//   **
                4'h8: data = 8'b00011000;	//   **
                4'h9: data = 8'b00011000;	//   **
                4'ha: data = 8'b11111000;	//*****
                4'hb: data = 8'b01111000;	// ****
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//    
                endcase
        end
        6'b001011: begin //K
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000110;	//**   **
                4'h3: data = 8'b11001100;	//**  **
                4'h4: data = 8'b11011000;	//** **
                4'h5: data = 8'b11110000;	//****
                4'h6: data = 8'b11100000;	//***
                4'h7: data = 8'b11100000;	//***
                4'h8: data = 8'b11110000;	//****
                4'h9: data = 8'b11011000;	//** **
                4'ha: data = 8'b11001100;	//**  **
                4'hb: data = 8'b11000110;	//**   **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//   
                endcase
        end
        6'b001100: begin //L
            case(row)
                4'h0: data = 8'b00000000;	    //
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000000;	//**
                4'h3: data = 8'b11000000;	//**
                4'h4: data = 8'b11000000;	//**
                4'h5: data = 8'b11000000;	//**
                4'h6: data = 8'b11000000;	//**
                4'h7: data = 8'b11000000;	//**
                4'h8: data = 8'b11000000;	//**
                4'h9: data = 8'b11000000;	//**
                4'ha: data = 8'b11111110;	//*******
                4'hb: data = 8'b11111110;	//*******
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b001101: begin //M
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000110;	//**   **
                4'h3: data = 8'b11000110;	//**   **
                4'h4: data = 8'b11101110;	//*** ***
                4'h5: data = 8'b11111110;	//*******
                4'h6: data = 8'b11010110;	//** * **
                4'h7: data = 8'b11000110;	//**   **
                4'h8: data = 8'b11000110;	//**   **
                4'h9: data = 8'b11000110;	//**   **
                4'ha: data = 8'b11000110;	//**   **
                4'hb: data = 8'b11000110;	//**   **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b001110: begin //N
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000110;	//**   **
                4'h3: data = 8'b11000110;	//**   **
                4'h4: data = 8'b11100110;	//***  **
                4'h5: data = 8'b11110110;	//**** **
                4'h6: data = 8'b11111110;	//*******
                4'h7: data = 8'b11011110;	//** ****
                4'h8: data = 8'b11001110;	//**  ***
                4'h9: data = 8'b11000110;	//**   **
                4'ha: data = 8'b11000110;	//**   **
                4'hb: data = 8'b11000110;	//**   **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
			endcase
        end  
        6'b001111: begin //O
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b01111100;	// *****
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **
                4'h6: data = 8'b11000110;	//**   **
                4'h7: data = 8'b11000110;	//**   **
                4'h8: data = 8'b11000110;	//**   **
                4'h9: data = 8'b11000110;	//**   **
                4'ha: data = 8'b11111110;	//*******
                4'hb: data = 8'b01111100;	// *****
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//  
                endcase
        end
        6'b010000: begin //P
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111100;	//******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **
                4'h6: data = 8'b11111110;	//*******
                4'h7: data = 8'b11111100;	//******   
                4'h8: data = 8'b11000000;	//**   
                4'h9: data = 8'b11000000;	//**   
                4'ha: data = 8'b11000000;	//**
                4'hb: data = 8'b11000000;	//**
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b010001: begin //Q
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111100;	// *****
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **
                4'h6: data = 8'b11000110;	//**   **
                4'h7: data = 8'b11000110;	//**   **  
                4'h8: data = 8'b11010110;	//** * **
                4'h9: data = 8'b11111110;	//*******
                4'ha: data = 8'b01101100;	// ** ** 
                4'hb: data = 8'b00000110;	//     **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b010010: begin //R
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111100;	//******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **
                4'h6: data = 8'b11111110;	//*******
                4'h7: data = 8'b11111100;	//******   
                4'h8: data = 8'b11011000;	//** **  
                4'h9: data = 8'b11001100;	//**  ** 
                4'ha: data = 8'b11000110;	//**   **
                4'hb: data = 8'b11000110;	//**   **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b010011: begin //S
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b01111100;	// *****
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b11000000;	//**   
                4'h5: data = 8'b11000000;	//**   
                4'h6: data = 8'b11111100;	//******
                4'h7: data = 8'b01111110;	// ******   
                4'h8: data = 8'b00000110;	//     **  
                4'h9: data = 8'b00000110;	//     **
                4'ha: data = 8'b11111110;	//*******  
                4'hb: data = 8'b01111100;	// ***** 
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end  
        6'b010100: begin //T
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111110;	//*******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b00110000;	//  **
                4'h5: data = 8'b00110000;	//  **
                4'h6: data = 8'b00110000;	//  **
                4'h7: data = 8'b00110000;	//  **   
                4'h8: data = 8'b00110000;	//  **  
                4'h9: data = 8'b00110000;	//  **
                4'ha: data = 8'b00110000;	//  **  
                4'hb: data = 8'b00110000;	//  **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b010101: begin //U
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000110;	//**   **
                4'h3: data = 8'b11000110;	//**   **
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **
                4'h6: data = 8'b11000110;	//**   **
                4'h7: data = 8'b11000110;	//**   **
                4'h8: data = 8'b11000110;	//**   **
                4'h9: data = 8'b11000110;	//**   **
                4'ha: data = 8'b11111110;	//*******
                4'hb: data = 8'b01111100;	// *****
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b010110: begin //V
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000110;	//**   **
                4'h3: data = 8'b11000110;	//**   **
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **
                4'h6: data = 8'b11000110;	//**   **
                4'h7: data = 8'b11000110;	//**   **
                4'h8: data = 8'b11000110;	//**   **
                4'h9: data = 8'b01101100;	// ** **
                4'ha: data = 8'b00111000;	//  ***  
                4'hb: data = 8'b00010000;	//   * 
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//   
                endcase
        end
        6'b010111: begin //W
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000110;	//**   **
                4'h3: data = 8'b11000110;	//**   **
                4'h4: data = 8'b11000110;	//**   **
                4'h5: data = 8'b11000110;	//**   **
                4'h6: data = 8'b11000110;	//**   **
                4'h7: data = 8'b11000110;	//**   **
                4'h8: data = 8'b11010110;	//** * **
                4'h9: data = 8'b11111110;	//*******
                4'ha: data = 8'b11101110;	//*** ***  
                4'hb: data = 8'b11000110;	//**   **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end  
        6'b011000: begin //X
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000110;	//**   **
                4'h3: data = 8'b11000110;	//**   **
                4'h4: data = 8'b01101100;	// ** ** 
                4'h5: data = 8'b00111000;	//  ***
                4'h6: data = 8'b00111000;	//  *** 
                4'h7: data = 8'b00111000;	//  ***
                4'h8: data = 8'b00111000;	//  ***
                4'h9: data = 8'b01101100;	// ** **
                4'ha: data = 8'b11000110;	//**   **  
                4'hb: data = 8'b11000110;	//**   **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	// 
                endcase
        end
        6'b011001: begin //Y
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11000110;	//**   **
                4'h3: data = 8'b11000110;	//**   **
                4'h4: data = 8'b01101100;	// ** ** 
                4'h5: data = 8'b00111000;	//  ***
                4'h6: data = 8'b00011000;	//   ** 
                4'h7: data = 8'b00011000;	//   **
                4'h8: data = 8'b00011000;	//   **
                4'h9: data = 8'b00011000;	//   **
                4'ha: data = 8'b00011000;	//   **  
                4'hb: data = 8'b00011000;	//   **
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b011010: begin //Z
            case(row)
                4'h0: data = 8'b00000000;	//
                4'h1: data = 8'b00000000;	//
                4'h2: data = 8'b11111110;	//*******
                4'h3: data = 8'b11111110;	//*******
                4'h4: data = 8'b00000110;	//     **  
                4'h5: data = 8'b00001100;	//    **
                4'h6: data = 8'b00011000;	//   ** 
                4'h7: data = 8'b00110000;	//  **
                4'h8: data = 8'b01100000;	// **
                4'h9: data = 8'b11000000;	//**
                4'ha: data = 8'b11111110;	//*******  
                4'hb: data = 8'b11111110;	//*******
                4'hc: data = 8'b00000000;	//
                4'hd: data = 8'b00000000;	//
                4'he: data = 8'b00000000;	//
                4'hf: data = 8'b00000000;	//
                endcase
        end
        6'b011011: begin //1
            case(row)
			4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b00011000;	//   **  
			4'h3: data = 8'b00111000;	//  ***
			4'h4: data = 8'b01111000;	// ****
			4'h5: data = 8'b00011000;	//   **
			4'h6: data = 8'b00011000;	//   **
			4'h7: data = 8'b00011000;	//   **
			4'h8: data = 8'b00011000;	//   **
			4'h9: data = 8'b00011000;	//   **
			4'ha: data = 8'b01111110;	// ******
			4'hb: data = 8'b01111110;	// ******
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
            endcase
        end
        6'b011100: begin //2
            case(row)
            4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b11111110;	//*******  
			4'h3: data = 8'b11111110;	//*******
			4'h4: data = 8'b00000110;	//     **
			4'h5: data = 8'b00000110;	//     **
			4'h6: data = 8'b11111110;	//*******
			4'h7: data = 8'b11111110;	//*******
			4'h8: data = 8'b11000000;	//**
			4'h9: data = 8'b11000000;	//**
			4'ha: data = 8'b11111110;	//*******
			4'hb: data = 8'b11111110;	//*******
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b011101: begin //3
            case(row)
            4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b11111110;	//*******  
			4'h3: data = 8'b11111110;	//*******
			4'h4: data = 8'b00000110;	//     **
			4'h5: data = 8'b00000110;	//     **
			4'h6: data = 8'b00111110;	//  *****
			4'h7: data = 8'b00111110;	//  *****
			4'h8: data = 8'b00000110;	//     **
			4'h9: data = 8'b00000110;	//     **
			4'ha: data = 8'b11111110;	//*******
			4'hb: data = 8'b11111110;	//*******
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b011110: begin //4
            case(row)
            4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b11000110;	//**   **  
			4'h3: data = 8'b11000110;	//**   **
			4'h4: data = 8'b11000110;	//**   **
			4'h5: data = 8'b11000110;	//**   **
			4'h6: data = 8'b11111110;	//*******
			4'h7: data = 8'b11111110;	//*******
			4'h8: data = 8'b00000110;	//     **
			4'h9: data = 8'b00000110;	//     **
			4'ha: data = 8'b00000110;	//     **
			4'hb: data = 8'b00000110;	//     **
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b011111: begin //5
            case(row)
            4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b11111110;	//*******  
			4'h3: data = 8'b11111110;	//*******
			4'h4: data = 8'b11000000;	//**
			4'h5: data = 8'b11000000;	//**
			4'h6: data = 8'b11111110;	//*******
			4'h7: data = 8'b11111110;	//*******
			4'h8: data = 8'b00000110;	//     **
			4'h9: data = 8'b00000110;	//     **
			4'ha: data = 8'b11111110;	//*******
			4'hb: data = 8'b11111110;	//*******
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b100000: begin //6
            case(row)
            4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b11111110;	//*******  
			4'h3: data = 8'b11111110;	//*******
			4'h4: data = 8'b11000000;	//**
			4'h5: data = 8'b11000000;	//**
			4'h6: data = 8'b11111110;	//*******
			4'h7: data = 8'b11111110;	//*******
			4'h8: data = 8'b11000110;	//**   **
			4'h9: data = 8'b11000110;	//**   **
			4'ha: data = 8'b11111110;	//*******
			4'hb: data = 8'b11111110;	//*******
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b100001: begin //7
            case(row)
            4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b11111110;	//*******  
			4'h3: data = 8'b11111110;	//*******
			4'h4: data = 8'b00000110;	//     **
			4'h5: data = 8'b00000110;	//     **
			4'h6: data = 8'b00000110;	//     **
			4'h7: data = 8'b00000110;	//     **
			4'h8: data = 8'b00000110;	//     **
			4'h9: data = 8'b00000110;	//     **
			4'ha: data = 8'b00000110;	//     **
			4'hb: data = 8'b00000110;	//     **
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b100010: begin //8
            case(row)
            4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b11111110;	//*******  
			4'h3: data = 8'b11111110;	//*******
			4'h4: data = 8'b11000110;	//**   **
			4'h5: data = 8'b11000110;	//**   **
			4'h6: data = 8'b11111110;	//*******
			4'h7: data = 8'b11111110;	//*******
			4'h8: data = 8'b11000110;	//**   **
			4'h9: data = 8'b11000110;	//**   **
			4'ha: data = 8'b11111110;	//*******
			4'hb: data = 8'b11111110;	//*******
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b100011: begin //9
            case(row)
            4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b11111110;	//*******  
			4'h3: data = 8'b11111110;	//*******
			4'h4: data = 8'b11000110;	//**   **
			4'h5: data = 8'b11000110;	//**   **
			4'h6: data = 8'b11111110;	//*******
			4'h7: data = 8'b11111110;	//*******
			4'h8: data = 8'b00000110;	//     **
			4'h9: data = 8'b00000110;	//     **
			4'ha: data = 8'b11111110;	//*******
			4'hb: data = 8'b11111110;	//*******
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
			endcase
        end
        6'b100100:begin //0
            case(row)
            4'h0: data = 8'b00000000;	//
			4'h1: data = 8'b00000000;	//
			4'h2: data = 8'b00111000;	//  ***  
			4'h3: data = 8'b01101100;	// ** **
			4'h4: data = 8'b11000110;	//**   **
			4'h5: data = 8'b11000110;	//**   **
			4'h6: data = 8'b11000110;	//**   **
			4'h7: data = 8'b11000110;	//**   **
			4'h8: data = 8'b11000110;	//**   **
			4'h9: data = 8'b11000110;	//**   **
			4'ha: data = 8'b01101100;	// ** **
			4'hb: data = 8'b00111000;	//  ***
			4'hc: data = 8'b00000000;	//
			4'hd: data = 8'b00000000;	//
			4'he: data = 8'b00000000;	//
			4'hf: data = 8'b00000000;	//
			endcase
	   end

        endcase
endmodule




